library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TPFINAL is
    Port ( ENVIAR : in  STD_LOGIC;
           MENSAJE : out  STD_LOGIC_VECTOR (11 downto 0));
end TPFINAL;

architecture Behavioral of TPFINAL is
--seniales

--

--declaracion componentes

--
begin


end Behavioral;

